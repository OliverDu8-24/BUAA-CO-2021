`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:17:09 10/22/2021
// Design Name:   splitter
// Module Name:   G:/MyWorkspace/Computer_Organization/ISE_Project/P0_L0_Splitter/splitter_tb.v
// Project Name:  P0_L0_Splitter
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: splitter
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module splitter_tb;

	// Inputs
	reg [31:0] A;

	// Outputs
	wire [7:0] O1;
	wire [7:0] O2;
	wire [7:0] O3;
	wire [7:0] O4;

	// Instantiate the Unit Under Test (UUT)
	splitter uut (
		.A(A), 
		.O1(O1), 
		.O2(O2), 
		.O3(O3), 
		.O4(O4)
	);

	initial begin
		// Initialize Inputs
		A = 32'b1000_0110_1101_1110_1111_0000_1010_0011;

		// Wait 100 ns for global reset to finish
		#5;
		$finish;
        
		// Add stimulus here

	end
      
endmodule

